LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;



ENTITY prom_a2l IS
	
	GENERIC
	(
		data_size		: INTEGER := 16;
		prom_size		: INTEGER := 256;
		addr_size		: INTEGER := 8
	);
	
	PORT
	(
		address		: IN STD_LOGIC_VECTOR(addr_size - 1 DOWNTO 0);
		
		data_out	: OUT STD_LOGIC_VECTOR(data_size - 1 DOWNTO 0)
	);
END prom_a2l;

--

ARCHITECTURE behavioral OF prom_a2l IS

	TYPE prom_memory IS ARRAY (0 TO prom_size - 1) OF STD_LOGIC_VECTOR(data_size - 1 DOWNTO 0);

	CONSTANT prom : prom_memory := 
	(
	"1110101010000000" ,
	"1110101110000000" ,
	"1110100010000000" ,
	"1110100110000000" ,
	"1110111010000000" ,
	"1110111110000000" ,
	"1110110010000000" ,
	"1110110110000000" ,
	"1110001010000000" ,
	"1110001110000000" ,
	"1110000010000000" ,
	"1110000110000000" ,
	"1110011010000000" ,
	"1110011110000000" ,
	"1110010010000000" ,
	"1110010110000000" ,
	"1111010101000000" ,
	"1111010111000000" ,
	"1111010001000000" ,
	"1111010011000000" ,
	"1111011101000000" ,
	"1111011111000000" ,
	"1111011001000000" ,
	"1111011011000000" ,
	"1111000101000000" ,
	"1111000111000000" ,
	"1111000001000000" ,
	"1111000011000000" ,
	"1111001101000000" ,
	"1111001111000000" ,
	"1111001001000000" ,
	"1111001011000000" ,
	"1010101000000000" ,
	"1010111000000000" ,
	"1010001000000000" ,
	"1010011000000000" ,
	"1011101000000000" ,
	"1011111000000000" ,
	"1011001000000000" ,
	"1011011000000000" ,
	"1000101000000000" ,
	"1000111000000000" ,
	"1000001000000000" ,
	"1000011000000000" ,
	"1001101000000000" ,
	"1001111000000000" ,
	"1001001000000000" ,
	"1001011000000000" ,
	"1101010100000000" ,
	"1101011100000000" ,
	"1101000100000000" ,
	"1101001100000000" ,
	"1101110100000000" ,
	"1101111100000000" ,
	"1101100100000000" ,
	"1101101100000000" ,
	"1100010100000000" ,
	"1100011100000000" ,
	"1100000100000000" ,
	"1100001100000000" ,
	"1100110100000000" ,
	"1100111100000000" ,
	"1100100100000000" ,
	"1100101100000000" ,
	"1111111010101000" ,
	"1111111010111000" ,
	"1111111010001000" ,
	"1111111010011000" ,
	"1111111011101000" ,
	"1111111011111000" ,
	"1111111011001000" ,
	"1111111011011000" ,
	"1111111000101000" ,
	"1111111000111000" ,
	"1111111000001000" ,
	"1111111000011000" ,
	"1111111001101000" ,
	"1111111001111000" ,
	"1111111001001000" ,
	"1111111001011000" ,
	"1111111110101000" ,
	"1111111110111000" ,
	"1111111110001000" ,
	"1111111110011000" ,
	"1111111111101000" ,
	"1111111111111000" ,
	"1111111111001000" ,
	"1111111111011000" ,
	"1111111100101000" ,
	"1111111100111000" ,
	"1111111100001000" ,
	"1111111100011000" ,
	"1111111101101000" ,
	"1111111101111000" ,
	"1111111101001000" ,
	"1111111101011000" ,
	"1111101010100000" ,
	"1111101011100000" ,
	"1111101000100000" ,
	"1111101001100000" ,
	"1111101110100000" ,
	"1111101111100000" ,
	"1111101100100000" ,
	"1111101101100000" ,
	"1111100010100000" ,
	"1111100011100000" ,
	"1111100000100000" ,
	"1111100001100000" ,
	"1111100110100000" ,
	"1111100111100000" ,
	"1111100100100000" ,
	"1111100101100000" ,
	"1111110101010000" ,
	"1111110101110000" ,
	"1111110100010000" ,
	"1111110100110000" ,
	"1111110111010000" ,
	"1111110111110000" ,
	"1111110110010000" ,
	"1111110110110000" ,
	"1111110001010000" ,
	"1111110001110000" ,
	"1111110000010000" ,
	"1111110000110000" ,
	"1111110011010000" ,
	"1111110011110000" ,
	"1111110010010000" ,
	"1111110010110000" ,
	"0001010110000000" ,
	"0001010010000000" ,
	"0001011110000000" ,
	"0001011010000000" ,
	"0001000110000000" ,
	"0001000010000000" ,
	"0001001110000000" ,
	"0001001010000000" ,
	"0001110110000000" ,
	"0001110010000000" ,
	"0001111110000000" ,
	"0001111010000000" ,
	"0001100110000000" ,
	"0001100010000000" ,
	"0001101110000000" ,
	"0001101010000000" ,
	"0000101011000000" ,
	"0000101001000000" ,
	"0000101111000000" ,
	"0000101101000000" ,
	"0000100011000000" ,
	"0000100001000000" ,
	"0000100111000000" ,
	"0000100101000000" ,
	"0000111011000000" ,
	"0000111001000000" ,
	"0000111111000000" ,
	"0000111101000000" ,
	"0000110011000000" ,
	"0000110001000000" ,
	"0000110111000000" ,
	"0000110101000000" ,
	"0101011000000000" ,
	"0101001000000000" ,
	"0101111000000000" ,
	"0101101000000000" ,
	"0100011000000000" ,
	"0100001000000000" ,
	"0100111000000000" ,
	"0100101000000000" ,
	"0111011000000000" ,
	"0111001000000000" ,
	"0111111000000000" ,
	"0111101000000000" ,
	"0110011000000000" ,
	"0110001000000000" ,
	"0110111000000000" ,
	"0110101000000000" ,
	"0010101100000000" ,
	"0010100100000000" ,
	"0010111100000000" ,
	"0010110100000000" ,
	"0010001100000000" ,
	"0010000100000000" ,
	"0010011100000000" ,
	"0010010100000000" ,
	"0011101100000000" ,
	"0011100100000000" ,
	"0011111100000000" ,
	"0011110100000000" ,
	"0011001100000000" ,
	"0011000100000000" ,
	"0011011100000000" ,
	"0011010100000000" ,
	"0000000101011000" ,
	"0000000101001000" ,
	"0000000101111000" ,
	"0000000101101000" ,
	"0000000100011000" ,
	"0000000100001000" ,
	"0000000100111000" ,
	"0000000100101000" ,
	"0000000111011000" ,
	"0000000111001000" ,
	"0000000111111000" ,
	"0000000111101000" ,
	"0000000110011000" ,
	"0000000110001000" ,
	"0000000110111000" ,
	"0000000110101000" ,
	"0000000001011000" ,
	"0000000001001000" ,
	"0000000001111000" ,
	"0000000001101000" ,
	"0000000000011000" ,
	"0000000000001000" ,
	"0000000000111000" ,
	"0000000000101000" ,
	"0000000011011000" ,
	"0000000011001000" ,
	"0000000011111000" ,
	"0000000011101000" ,
	"0000000010011000" ,
	"0000000010001000" ,
	"0000000010111000" ,
	"0000000010101000" ,
	"0000010101100000" ,
	"0000010100100000" ,
	"0000010111100000" ,
	"0000010110100000" ,
	"0000010001100000" ,
	"0000010000100000" ,
	"0000010011100000" ,
	"0000010010100000" ,
	"0000011101100000" ,
	"0000011100100000" ,
	"0000011111100000" ,
	"0000011110100000" ,
	"0000011001100000" ,
	"0000011000100000" ,
	"0000011011100000" ,
	"0000011010100000" ,
	"0000001010110000" ,
	"0000001010010000" ,
	"0000001011110000" ,
	"0000001011010000" ,
	"0000001000110000" ,
	"0000001000010000" ,
	"0000001001110000" ,
	"0000001001010000" ,
	"0000001110110000" ,
	"0000001110010000" ,
	"0000001111110000" ,
	"0000001111010000" ,
	"0000001100110000" ,
	"0000001100010000" ,
	"0000001101110000" ,
	"0000001101010000" 
	);

BEGIN
	data_out <= prom(CONV_INTEGER(address));
	
END behavioral;

